library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity DECODER2_4 is 
	Port( 
			S: in STD_LOGIC_VECTOR(1 downto 0);
			Y:	 out STD_LOGIC_VECTOR(3 downto 0));
end DECODER2_4;


architecture Behavioral of DECODER2_4 is

begin
	process (S)
    begin
        case S is
            when "00" =>
                Y <= "1101";
            when "01" =>
                Y <= "1011";
            when "10" =>
                Y <= "0111";
            when "11" =>
                Y <= "1110";
				when others =>
                Y <= "1111"; 
        end case;
   end process;
	  
end Behavioral;