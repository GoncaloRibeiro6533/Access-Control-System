library IEEE;
use IEEE.std_logic_1164.all;

entity SLCDC_TB is
end SLCDC_TB;

architecture testbench of SLCDC_TB is
    -- Component declarations
    component SLCDC is
        port (
            MCLK, reset : in std_logic;
            NOT_SS, SCLK, SDX : in std_logic;
            WrL : out std_logic;
            Dout : out std_logic_vector(4 downto 0)
        );
    end component;

    -- Signal declarations
    signal MCLK_in, reset_in, NOT_SS_in, SCLK_in, SDX_in : std_logic;
    signal WrL_out : std_logic;
    signal Dout_out : std_logic_vector(4 downto 0);

begin
    -- Instantiate the SLCDC
    UUT: SLCDC port map (
        MCLK => MCLK_in,
        reset => reset_in,
        NOT_SS => NOT_SS_in,
        SCLK => SCLK_in,
        SDX => SDX_in,
        WrL => WrL_out,
        Dout => Dout_out
    );

    -- Stimulus process
    stimulus: process
    begin
        -- Initialize signals
        MCLK_in <= '0';
        reset_in <= '1';
        NOT_SS_in <= '0';
        SCLK_in <= '0';
        SDX_in <= '0';
        wait for 10 ns;

        -- Release reset
        reset_in <= '0';
        wait for 10 ns;

        -- Apply stimuli
        NOT_SS_in <= '1';
        SCLK_in <= '1';
        SDX_in <= '1';
        wait for 10 ns;

        -- End the simulation
        wait;
    end process;

 

end testbench;
