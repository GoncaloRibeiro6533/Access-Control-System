library IEEE;
use IEEE.std_logic_1164.all;

entity DoorController_TB is
end DoorController_TB;

architecture testbench of DoorController_TB is
    -- Component declarations
    component DoorController is
        port (
            Dval, clk, reset, Sclose, Sopen, Psensor : in std_logic;
            OnOff, done, OpenClose : out std_logic;
            Din : in std_logic_vector (4 downto 0);
            Dout : out std_logic_vector (4 downto 0)
        );
    end component;

    -- Signal declarations
    signal Dval_in, clk_in, reset_in, Sclose_in, Sopen_in, Psensor_in : std_logic;
    signal OnOff_out, done_out, OpenClose_out : std_logic;
    signal Din_in : std_logic_vector (4 downto 0);
    signal Dout_out : std_logic_vector (4 downto 0);

begin
    -- Instantiate the DoorController
    UUT: DoorController port map (
        Dval => Dval_in,
        clk => clk_in,
        reset => reset_in,
        Sclose => Sclose_in,
        Sopen => Sopen_in,
        Psensor => Psensor_in,
        OnOff => OnOff_out,
        done => done_out,
        OpenClose => OpenClose_out,
        Din => Din_in,
        Dout => Dout_out
    );

    -- Stimulus process
    stimulus: process
    begin
        -- Initialize signals
        Dval_in <= '0';
        clk_in <= '0';
        reset_in <= '1';
        Sclose_in <= '0';
        Sopen_in <= '0';
        Psensor_in <= '0';
        Din_in <= (others => '0');
        wait for 10 ns;

        -- Release reset
        reset_in <= '0';
        wait for 10 ns;

        -- Apply stimuli
        Dval_in <= '1';
        clk_in <= '1';
        wait for 10 ns;

        Sclose_in <= '1';
        wait for 10 ns;

        Sopen_in <= '1';
        Din_in <= "00001";
        wait for 10 ns;

        Psensor_in <= '1';
        wait for 10 ns;

        Sclose_in <= '0';
        wait for 10 ns;

        Psensor_in <= '0';
        wait for 10 ns;

        Sopen_in <= '0';
        Din_in <= "00000";
        wait for 10 ns;

        Dval_in <= '0';
        wait for 10 ns;
	end process;

end testbench;
